`define CPU_ARCH 32
module pc_add(
		input [`CPU_ARCH -1:0] pc,
		output [`CPU_ARCH-1:0] pc_next); 
	
	assign pc_next = pc+4;
		
endmodule 
