

module core(
		input clk_i,
		input rst_i,
		input 
